module andstr(x,y,z);
input x,y;
output z;
and gl(z,x,y);
endmodule
