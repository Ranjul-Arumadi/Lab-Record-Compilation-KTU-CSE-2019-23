module andstr(x,y,z);
input x,y;
output z;
or gl(z,x,y);
endmodule
